`timescale 1ns / 1ps

module InsMEM(
        input [31:0] curPC,      //PC值
        output reg[7:0] op,      //操作码位段
        output reg[2:0] funct3,  //3位功能码位段
        output reg[6:0] funct7,  //7位功能码位段
        output reg[4:0] rs1,     //rs1地址位段
        output reg[4:0] rs2,     //rs2地址位段
        output reg[4:0] rd,      //rd地址位段
        output reg[24:0] imm,    //立即数位段传给extend模块拼接扩展
        output reg [31:0] instr  //读取得到32位指令
    );
    reg [7:0] rom[128:0];  //存储器定义必须用reg类型，存储器存储单元8位长度，共128个存储单元，可以存32条指令

    // 加载数据到存储器rom
    initial begin
        //$readmemb("X://rom.txt", rom);
        {rom[3],rom[2],rom[1],rom[0]}     = 32'b00000000100000000000000010010011;
        {rom[7],rom[6],rom[5],rom[4]}     = 32'b00000000001000000110000100010011;
        {rom[11],rom[10],rom[9],rom[8]}   = 32'b00000000000100010000000110110011;
        {rom[15],rom[14],rom[13],rom[12]} = 32'b01000000001000011000001010110011;
        {rom[19],rom[18],rom[17],rom[16]} = 32'b00000000001000101111001000110011;
        {rom[23],rom[22],rom[21],rom[20]} = 32'b00000000001000100110010000110011;
        {rom[27],rom[26],rom[25],rom[24]} = 32'b00000000000101000001010000010011;
        {rom[31],rom[30],rom[29],rom[28]} = 32'b11111110000101000001111011100011;
        {rom[35],rom[34],rom[33],rom[32]} = 32'b00000000010000010010001100010011;
        {rom[39],rom[38],rom[37],rom[36]} = 32'b00000000000000110010001110010011;
        {rom[43],rom[42],rom[41],rom[40]} = 32'b00000000100000111000001110010011;
        {rom[47],rom[46],rom[45],rom[44]} = 32'b11111110000100111000111011100011;
        {rom[51],rom[50],rom[49],rom[48]} = 32'b00000000001000001010001000100011;
        {rom[55],rom[54],rom[53],rom[52]} = 32'b00000000010000001010010010000011;
        {rom[59],rom[58],rom[57],rom[56]} = 32'b11111111111000000000010100010011;
        {rom[63],rom[62],rom[61],rom[60]} = 32'b00000000000101010000010100010011;
        {rom[67],rom[66],rom[65],rom[64]} = 32'b11111110000001010100111011100011;
        {rom[71],rom[70],rom[69],rom[68]} = 32'b00000000001000010111010110010011;
        {rom[75],rom[74],rom[73],rom[72]} = 32'b00000000100000000000010001101111;
        {rom[79],rom[78],rom[77],rom[76]} = 32'b00000000100000000000010001101111;
        {rom[83],rom[82],rom[81],rom[80]} = 32'b00000000000000000000000001100011;

        op = 7'b0000000;
        funct3 = 3'b000;
        funct7 = 7'b0000000;
        rs1 = 5'b00000;
        rs2 = 5'b00000;
        imm = 20'b00000000000000000000;
    end

    //小端模式,PC改变就取指令
    always@(curPC)
    begin
        //取指令
        begin
            instr[7:0] = rom[curPC];
            instr[15:8] = rom[curPC + 1];
            instr[23:16] = rom[curPC + 2];
            instr[31:24] = rom[curPC + 3];
        end 
    end
    //切割指令
    always@(instr) 
    begin
        op = instr[6:0];
        rs1 = instr[19:15];
        rs2 = instr[24:20];
        rd = instr[11:7];
        funct3 = instr[14:12];
        funct7 = instr[31:26];
        imm = instr[31:7];
    end

endmodule